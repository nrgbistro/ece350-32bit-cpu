module not_equal(
    output out,
    input [31:0] a, b);


endmodule
