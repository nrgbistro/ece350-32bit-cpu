module multControl(
    output [1:0] productInputCode,
    output sub,
    input [2:0] opCode,
    input count0bool);

endmodule
