module regfile (
	clock,
	ctrl_writeEnable, ctrl_reset, ctrl_writeReg,
	ctrl_readRegA, ctrl_readRegB, data_writeReg,
	data_readRegA, data_readRegB);

	input clock, ctrl_writeEnable, ctrl_reset;
	input [4:0] ctrl_writeReg, ctrl_readRegA, ctrl_readRegB;
	input [31:0] data_writeReg;
	output [31:0] data_readRegA, data_readRegB;

    // 32bit register selection bus for each 1bit register
    wire [31:0][31:0] regOut;
    wire [31:0] triStateSelectA, triStateSelectB, selectWriteRegDecoded;

    decoder32 decoderA(triStateSelectA, 1'b1, ctrl_readRegA);
    decoder32 decoderB(triStateSelectB, 1'b1, ctrl_readRegB);
    decoder32 selectWriteReg(selectWriteRegDecoded, ctrl_writeEnable, ctrl_writeReg);

    genvar i;
    for (i = 0; i < 32; i = i + 1) begin : registers
        // Don't allow reg0 to be written to
        if(i == 0) begin
            register32 reg32(regOut[i], data_writeReg, clock, 1'b0, ctrl_reset);
        end else begin
            register32 reg32(regOut[i], data_writeReg, clock, selectWriteRegDecoded[i], ctrl_reset);
        end
        tri_state32 triStateA(data_readRegA, triStateSelectA[i], regOut[i]);
        tri_state32 triStateB(data_readRegB, triStateSelectB[i], regOut[i]);
    end

endmodule
