module resetDetection(
    output rst,
    input div, mult, clock);


endmodule
