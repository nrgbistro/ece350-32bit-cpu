module cla_32(
    output [3:0] carry,
    input [3:0] PG, GG);


    assign carry[0] = 0;

endmodule
