module cla
    (output [31:0] sum,
    input [31:0] a, b);

endmodule
