module adder_8(
    output Cout, PG, GG,
    input [7:0] a, b,
    input Cin);

endmodule
