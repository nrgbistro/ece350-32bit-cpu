module processorControl(
    output o1,
    input [5:0] opCode);

endmodule
