module resetDetection(
    output rst,
    input div, mult, clock);

    assign rst = 1'b0;

endmodule
