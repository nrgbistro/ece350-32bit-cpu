module cla(
    output [31:0] Cout, Cin,
    input [31:0] a, b, p, g);

endmodule
