module Timer(
    output reg [31:0] t,
    input clock, reset)


endmodule
